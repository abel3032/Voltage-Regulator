** Profile: "SCHEMATIC1-ripl"  [ d:\proiectul_meu\proiect-PSpiceFiles\SCHEMATIC1\ripl.sim ] 

** Creating circuit file "ripl.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Profile Libraries :
* Local Libraries :
.LIB "C:/Users/alber/OneDrive/Desktop/librarii_proiect/Lib_ModelePSpice_Anexa_1/Modele_A1_lib/SMLS14BET.lib" 
.LIB "C:/Users/alber/OneDrive/Desktop/librarii_proiect/Lib_ModelePSpice_Anexa_1/Modele_A1_lib/BC856B.lib" 
.LIB "C:/Users/alber/OneDrive/Desktop/librarii_proiect/Lib_ModelePSpice_Anexa_1/Modele_A1_lib/BZX84C5V6.lib" 
.LIB "C:/Users/alber/OneDrive/Desktop/librarii_proiect/Lib_ModelePSpice_Anexa_1/Modele_A1_lib/BC846B.lib" 
.LIB "C:/Users/alber/OneDrive/Desktop/librarii_proiect/Lib_ModelePSpice_Anexa_1/Modele_A1_lib/MJD31CG.lib" 
.LIB "C:/Users/alber/OneDrive/Desktop/librarii_proiect/Lib_ModelePSpice_Anexa_1/Modele_A1_lib/BC817-25.lib" 
.LIB "C:/Users/alber/OneDrive/Desktop/librarii_proiect/Lib_ModelePSpice_Anexa_1/Modele_A1_lib/BZX84C2V7.lib" 
.LIB "C:/Users/alber/OneDrive/Desktop/librarii_proiect/Lib_ModelePSpice_Anexa_1/Modele_A1_lib/BZX84C5V1.lib" 
.LIB "C:/Users/alber/OneDrive/Desktop/librarii_proiect/Lib_ModelePSpice_Anexa_1/Modele_A1_lib/BZX84C6V8.lib" 
* From [PSPICE NETLIST] section of C:\Users\alber\AppData\Roaming\SPB_Data\cdssetup\OrCAD_PSpice/16.6.0/PSpice.ini file:
.lib "nomd.lib" 

*Analysis directives: 
.TRAN  0 5ms 0 
.OPTIONS ADVCONV
.PROBE64 V(alias(*)) I(alias(*)) W(alias(*)) D(alias(*)) NOISE(alias(*)) 
.INC "..\SCHEMATIC1.net" 


.END
